`timescale 1ns/1ps

module Max_Data_tb();
	parameter t = 10;
	parameter data_width = 32;
	parameter R = 2;
	parameter C = 2;

	reg[data_width*R*C:0] In;
	wire[data_width-1:0] max_data;

	initial begin
		#t In = 'b0011_1111_1100_0000_0000_0000_0000_0000_0100_0000_0000_0000_0000_0000_0000_0000_0100_0000_0010_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
		#(t*2) In = 'b0011_1110_0000_0010_0000_1100_0100_1010_0100_0001_0010_0110_0110_0110_0110_0110_0100_0000_1111_1001_1001_1001_1001_1010_0011_1101_1110_0011_0101_0011_1111_1000;
		#(t*4) $finish;
	end

	Max_Data #(data_width, R, C) DUT(max_data, In);

endmodule

/*
In = [1.5 2 2.5 0]
=> max_data = 'b0100_0000_0010_0000_0000_0000_0000_0000 (2.5)
In = [0.127 10.4 7.8 0.111]
=> max_data = 'b0100_0001_0010_0110_0110_0110_0110_0110
*/
